module bin_to_sseg (
  // input wire CLOCK,
  input wire [3:0] BIN,
  output wire [6:0] HEX
);

assign HEX = 
  (BIN == 4'b0000) ? 7'b1000000 :
  (BIN == 4'b0001) ? 7'b1111001 :
  (BIN == 4'b0010) ? 7'b0100100 :
  (BIN == 4'b0011) ? 7'b0110000 :
  (BIN == 4'b0100) ? 7'b0011001 :
  (BIN == 4'b0101) ? 7'b0010010 :
  (BIN == 4'b0110) ? 7'b0000010 :
  (BIN == 4'b0111) ? 7'b1111000 :
  (BIN == 4'b1000) ? 7'b0000000 :
  (BIN == 4'b1001) ? 7'b0010000 :
  (BIN == 4'b1010) ? 7'b0001000 :
  (BIN == 4'b1011) ? 7'b0000011 :
  (BIN == 4'b1100) ? 7'b1000110 :
  (BIN == 4'b1101) ? 7'b0100001 :
  (BIN == 4'b1110) ? 7'b0000110 : 7'b0001110;
  // (BIN == 4'b1111) ? 7'b0001110 : 7'b0101011;

endmodule
