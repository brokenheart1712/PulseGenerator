module bin_to_sseg (
  // input wire CLOCK,
  input wire [3:0] BIN,
  output wire [6:0] HEX
);

assign HEX = 
  (BIN == 4'b0000) ? 7'b1000000 : // 0
  (BIN == 4'b0001) ? 7'b1111001 : // 1
  (BIN == 4'b0010) ? 7'b0100100 : // 2
  (BIN == 4'b0011) ? 7'b0110000 : // 3
  (BIN == 4'b0100) ? 7'b0011001 : // 4
  (BIN == 4'b0101) ? 7'b0010010 : // 5
  (BIN == 4'b0110) ? 7'b0000010 : // 6
  (BIN == 4'b0111) ? 7'b1111000 : // 7
  (BIN == 4'b1000) ? 7'b0000000 : // 8
  (BIN == 4'b1001) ? 7'b0010000 : // 9
  (BIN == 4'b1010) ? 7'b1001000 : // n
  (BIN == 4'b1011) ? 7'b0000011 : // b
  (BIN == 4'b1100) ? 7'b1000110 : // c
  (BIN == 4'b1101) ? 7'b0100001 : // d
  (BIN == 4'b1110) ? 7'b0000110 : // e
                     7'b1111111;  // off

endmodule
